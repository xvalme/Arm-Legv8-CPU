module gates();

wire out0, out1, out2;
reg in1, in2, in3;

initial begin